/* datatypes.sv
 */

